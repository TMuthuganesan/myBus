`timescale 1ns/1ps
package myPkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  `include "transactionBaseClasses.sv"
  `include "transactions.sv"
  `include "sequencer.sv"
  `include "driver.sv"
  `include "monitor.sv"
  `include "scoreboard.sv"
  `include "agent.sv"
  `include "env.sv"
  `include "cpuWrSeq.sv"
  `include "directedCpuWrSeq.sv"
  `include "cpuRdSeq.sv"
  `include "baseTest.sv"
  `include "cpuWrTest.sv"
  `include "cpuRdTest.sv"
  `include "cpuWrRdTest.sv"
  `include "directedCpuWrTest.sv"
endpackage
